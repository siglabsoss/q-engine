// address decoder for the permutation network
// consumes destination address and produces source address

module perm_full_addr_dat_1_1 (
    input  [67:0] t_0_dat,
    output [67:0] i_0_dat,
    input clk, reset_n
);

assign i_0_dat = t_0_dat;

endmodule
