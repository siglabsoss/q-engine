

module cfg_ctrl_ (


    input clk, reset_n
);

endmodule
